module exe(

);


endmodule
